module dummy (/*AUTOARG*/);
            /*AUTOINPUT*/
            /*AUTOOUTPUT*/
            /*AUTOWIRE*/
            /*AUTOREG*/
endmodule